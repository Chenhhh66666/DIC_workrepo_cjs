`define WIDTH 32
`define DEPTH 9  //2的9次方=512
`define PATTERN "Standard"  //Standard,FWFT两种模式
`define THRESHOLD 10   //设置水位
`define FIFO_CNT_MAX 511