`define WIDTH 32
`define DEPTH 9  //2的9次方=512
`define PATTERN "Standard"  //Standard,FWFT两种模式
`define FIFO_CNT_MAX 511
`define full_threshold 500
`define empty_threshold 20