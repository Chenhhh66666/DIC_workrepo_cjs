`define DEPTH 3072 //���
`define ADDR 12  //��Ӧλ���ַ����
`define WIDTH 32  //����λ��
`define CLASH "WRITEFIRST"  //��ͻģʽ��NOCHANEG,READ,WRITE
`define CLASHB "READFIRST"  //��ͻģʽ��NOCHANEG,READ,WRITE
`define RAM_STYLE "block"
//`define WAVETYPE "TRI"  //TRI���ǲ� SIN���Ҳ� SQU����
