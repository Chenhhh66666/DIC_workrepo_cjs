`define DEPTH 1024 //深度
`define ADDR 10  //1024对应10位宽地址输入
`define WIDTH 32  //数据位宽
`define CLASH "NOCHANGE"  //冲突模式。NOCHANEG,READFIRST,WRITEFIRST
