parameter DEPTH = 1024;
parameter ADDR = 10;  //10位宽地址数，对应1024个地址
parameter WIDTH = 32;